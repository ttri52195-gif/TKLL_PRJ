/* verilator lint_off MULTITOP */

`timescale 1ns / 1ns

module Shift_Left_2(
    input [31:0] inp,
    output [31:0] out
);

    assign out = (inp << 2);
    
endmodule
